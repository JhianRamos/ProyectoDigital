module interfaz(msg,
					  Mostrar_10,
					  Mostrar_11,
					  Mostrar_12,
					  Mostrar_13,
					  Mostrar_14,
					  Mostrar_15,
					  Mostrar_16,
					  Mostrar_17,
					  Mostrar_18,
					  Mostrar_19,
					  Mostrar_110,
					  Mostrar_111,
					  Mostrar_112,
					  Mostrar_113,
					  Mostrar_114,
					  Mostrar_115,
					  Mostrar_20,
					  Mostrar_21,
					  Mostrar_22,
					  Mostrar_23,
					  Mostrar_24,
					  Mostrar_25,
					  Mostrar_26,
					  Mostrar_27,
					  Mostrar_28,
					  Mostrar_29,
					  Mostrar_210,
					  Mostrar_211,
					  Mostrar_212,
					  Mostrar_213,
					  Mostrar_214,
					  Mostrar_215);
	

    input [4:0]msg;
    output reg [8:0] Mostrar_10;
    output reg [8:0] Mostrar_11;
    output reg [8:0] Mostrar_12;
    output reg [8:0] Mostrar_13;
    output reg [8:0] Mostrar_14;
    output reg [8:0] Mostrar_15;
    output reg [8:0] Mostrar_16;
    output reg [8:0] Mostrar_17;
    output reg [8:0] Mostrar_18;
    output reg [8:0] Mostrar_19;
    output reg [8:0] Mostrar_110;
    output reg [8:0] Mostrar_111;
    output reg [8:0] Mostrar_112;
    output reg [8:0] Mostrar_113;
    output reg [8:0] Mostrar_114;
    output reg [8:0] Mostrar_115;
    output reg [8:0] Mostrar_20;
    output reg [8:0] Mostrar_21;
    output reg [8:0] Mostrar_22;
    output reg [8:0] Mostrar_23;
    output reg [8:0] Mostrar_24;
    output reg [8:0] Mostrar_25;
    output reg [8:0] Mostrar_26;
    output reg [8:0] Mostrar_27;
    output reg [8:0] Mostrar_28;
    output reg [8:0] Mostrar_29;
    output reg [8:0] Mostrar_210;
    output reg [8:0] Mostrar_211;
    output reg [8:0] Mostrar_212;
    output reg [8:0] Mostrar_213;
    output reg [8:0] Mostrar_214;
    output reg [8:0] Mostrar_215;


always
 begin

					  Mostrar_10=9'h120; //es
					  Mostrar_11=9'h141; //A
					  Mostrar_12=9'h13A; //:
					  Mostrar_13=9'h150; //P
					  Mostrar_14=9'h172; //r
					  Mostrar_15=9'h16F; //o
					  Mostrar_16=9'h167; //g
					  Mostrar_17=9'h172; //r
					  Mostrar_18=9'h161; //a
					  Mostrar_19=9'h16D;//m
					  Mostrar_110=9'h161; //a
					  Mostrar_111=9'h172; //r
					  Mostrar_112=9'h120;//es
					  Mostrar_113=9'h120;//es
					  Mostrar_114=9'h120;//es
					  Mostrar_115=9'h120;//es
					  Mostrar_20=9'h142;//B
					  Mostrar_21=9'h13A;//:
					  Mostrar_22=9'h152;//R
					  Mostrar_23=9'h165;//e
					  Mostrar_24=9'h169;//i
					  Mostrar_25=9'h16E;//n
					  Mostrar_26=9'h169;//i
					  Mostrar_27=9'h163;//c
					  Mostrar_28=9'h169;//i
					  Mostrar_29=9'h161;//a
					  Mostrar_210=9'h172;//r
					  Mostrar_211=9'h120;
					  Mostrar_212=9'h120;
					  Mostrar_213=9'h120;
					  Mostrar_214=9'h120;
					  Mostrar_215=9'h120;
				
					
//if (msg==4'hB) begin
//					  Mostrar_10=9'h120; //es
//					  Mostrar_11=9'h147; //G
//					  Mostrar_12=9'h161; //a
//					  Mostrar_13=9'h174; //t
//					  Mostrar_14=9'h16F; //o
//					  Mostrar_15=9'h120; //es
//					  Mostrar_16=9'h131; //1
//					  Mostrar_17=9'h12E; //.
//					  Mostrar_18=9'h120; //es
//					  Mostrar_19=9'h170; //P
//					  Mostrar_110=9'h165; //e
//					  Mostrar_111=9'h173; //s
//					  Mostrar_112=9'h16F;//o
//					  Mostrar_113=9'h120;//es
//					  Mostrar_114=9'h120;//es
//					  Mostrar_115=9'h120;//es
//					  Mostrar_20=9'h165;//e
//					  Mostrar_21=9'h16E;//n
//					  Mostrar_22=9'h120;//es
//					  Mostrar_23=9'h16B;//k
//					  Mostrar_24=9'h167;//g
//					  Mostrar_25=9'h12E;//.
//					  Mostrar_26=9'h120;
//					  Mostrar_27=9'h120;
//					  Mostrar_28=9'h120;
//					  Mostrar_29=9'h120;
//					  Mostrar_210=9'h120;
//					  Mostrar_211=9'h120;
//					  Mostrar_212=9'h120;
//					  Mostrar_213=9'h120;
//					  Mostrar_214=9'h120;
//					  Mostrar_215=9'h120;
//					end
		end

endmodule
